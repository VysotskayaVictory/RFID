`define CMD_NONE 0
`define CMD_START 1
`define CMD_A 2
`define CMD_FIN_A 3 
`define CMD_M 4 
`define CMD_FIN 5
`define WIDTH 64
`define KEY_WIDTH 256
`define LEN_WIDTH 64
`define BYTE_SIZE 8
`define STATE_WIDTH 5