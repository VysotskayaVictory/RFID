`define CMD_NONE 0
`define CMD_START_A 1
`define CMD_A 2
`define CMD_FIN_A 3
`define CMD_START_M 4 
`define CMD_DOUBLE_M 5
`define CMD_FIN_M 6
`define CMD_FIN 7
`define WIDTH 64
`define LOG_WIDTH 6
`define KEY_WIDTH 256
`define LEN_WIDTH 32
`define BYTE_SIZE 8 
`define STATE_WIDTH 7



